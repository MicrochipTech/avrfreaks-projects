// megafunction wizard: %LPM_LATCH%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_latch 

// ============================================================
// File Name: lpm_latch0.v
// Megafunction Name(s):
// 			lpm_latch
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 6.1 Build 201 11/27/2006 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2006 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module lpm_latch0 (
	data,
	gate,
	q);

	input	[8:0]  data;
	input	  gate;
	output	[8:0]  q;

	wire [8:0] sub_wire0;
	wire [8:0] q = sub_wire0[8:0];

	lpm_latch	lpm_latch_component (
				.data (data),
				.gate (gate),
				.q (sub_wire0),
				.aclr (1'b0),
				.aconst (1'b0),
				.aset (1'b0));
	defparam
		lpm_latch_component.lpm_type = "LPM_LATCH",
		lpm_latch_component.lpm_width = 9;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: aset NUMERIC "0"
// Retrieval info: PRIVATE: nBit NUMERIC "9"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_LATCH"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "9"
// Retrieval info: USED_PORT: data 0 0 9 0 INPUT NODEFVAL data[8..0]
// Retrieval info: USED_PORT: gate 0 0 0 0 INPUT NODEFVAL gate
// Retrieval info: USED_PORT: q 0 0 9 0 OUTPUT NODEFVAL q[8..0]
// Retrieval info: CONNECT: @data 0 0 9 0 data 0 0 9 0
// Retrieval info: CONNECT: q 0 0 9 0 @q 0 0 9 0
// Retrieval info: CONNECT: @gate 0 0 0 0 gate 0 0 0 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch0.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch0.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch0.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch0.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch0_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch0_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
